module findSign(output sign,input s1,input s2);
    assign sign = s1^s2;
endmodule