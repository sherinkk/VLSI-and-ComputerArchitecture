`include "adder.v"
module top;

reg [31:0] a,b;
wire [31:0] out;


adder s_1 (a,b,out);

initial 
begin
    a = 32'b01000000101000000000000000000000; //5
    b = 32'b01000001000000000000000000000000; //8
    #10 b=32'b11000000010000000000000000000000;//-3
    #10 b=32'b11000001000000000000000000000000;//-8
    #10 b=32'b11000001001000000000000000000000;//-10
    #10 b=32'b11000001000100000000000000000000;//-9
        a=32'b01000001000100000000000000000000;//+9
    #10 a=32'b01111111100000000000000000000000;
        b=32'b01011100101000000000000000000000;
    #10 a=32'b01000001010100000000000000000000;
        b=32'b01000000010000000000000000000000;
        



end

initial
    $monitor($time," a = %b; b = %b; out = %b;",a,b,out);
endmodule
