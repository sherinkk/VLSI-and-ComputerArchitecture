`include "WM.v"
module top;

	reg [31:0] a,b;
	wire[64:0]f_sum;
	
	WM wm1(a,b,f_sum);
	initial 
		begin
			a=32'b00000000000000000000010000000000;
			b=32'b00000000000000000000000000000001;
			#10 a=32'b00000000000000000000100000000011;
			#10 a=32'b00000000000000000000100000000010;
			#10 b=32'b00000000000000000000000000000010;
			#10 b=32'b00000000000000000000000000000011;
			/*#10 b=8'b00000011;
			#10 a=8'b10000001;
				b=8'b00000111;*/
		end
	
	initial
		begin
			$monitor("%b x %b  = %d", a, b,f_sum);
		end
		
endmodule
